module dut(
	input [17:0] a,
	output [17:0] z
);
	assign z = a;
endmodule
